UFM_NONE_inst : UFM_NONE PORT MAP (
		arclk	 => arclk_sig,
		ardin	 => ardin_sig,
		arshft	 => arshft_sig,
		drclk	 => drclk_sig,
		drdin	 => drdin_sig,
		drshft	 => drshft_sig,
		erase	 => erase_sig,
		oscena	 => oscena_sig,
		program	 => program_sig,
		busy	 => busy_sig,
		drdout	 => drdout_sig,
		osc	 => osc_sig,
		rtpbusy	 => rtpbusy_sig
	);
